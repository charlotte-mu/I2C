module lcd_rom(
	input [9:0] address,
	output [7:0] data_out
);
reg [7:0]rom[1023:0];
assign data_out = rom[address];
initial
begin
		rom[0]   	<= 8'hff;
		rom[1]   	<= 8'hff;
		rom[2]   	<= 8'hff;
		rom[3]   	<= 8'hff;
		rom[4]   	<= 8'hff;
		rom[5]   	<= 8'hff;
		rom[6]   	<= 8'hff;
		rom[7]   	<= 8'hff;
		rom[8]   	<= 8'hff;
		rom[9]   	<= 8'hff;
		rom[10]   	<= 8'hff;
		rom[11]   	<= 8'hff;
		rom[12]   	<= 8'hff;
		rom[13]   	<= 8'hff;
		rom[14]   	<= 8'hff;
		rom[15]   	<= 8'hff;
		rom[16]   	<= 8'hff;
		rom[17]   	<= 8'hff;
		rom[18]   	<= 8'hff;
		rom[19]   	<= 8'hff;
		rom[20]   	<= 8'hff;
		rom[21]   	<= 8'hff;
		rom[22]   	<= 8'hff;
		rom[23]   	<= 8'hff;
		rom[24]   	<= 8'hff;
		rom[25]   	<= 8'hff;
		rom[26]   	<= 8'hff;
		rom[27]   	<= 8'hff;
		rom[28]   	<= 8'hff;
		rom[29]   	<= 8'hff;
		rom[30]   	<= 8'hff;
		rom[31]   	<= 8'hff;
		rom[32]   	<= 8'hff;
		rom[33]   	<= 8'hff;
		rom[34]   	<= 8'hff;
		rom[35]   	<= 8'hff;
		rom[36]   	<= 8'hff;
		rom[37]   	<= 8'hff;
		rom[38]   	<= 8'hff;
		rom[39]   	<= 8'hff;
		rom[40]   	<= 8'hff;
		rom[41]   	<= 8'hff;
		rom[42]   	<= 8'hff;
		rom[43]   	<= 8'hff;
		rom[44]   	<= 8'hff;
		rom[45]   	<= 8'hff;
		rom[46]   	<= 8'hff;
		rom[47]   	<= 8'hff;
		rom[48]   	<= 8'hff;
		rom[49]   	<= 8'hff;
		rom[50]   	<= 8'hff;
		rom[51]   	<= 8'hff;
		rom[52]   	<= 8'hff;
		rom[53]   	<= 8'hff;
		rom[54]   	<= 8'hff;
		rom[55]   	<= 8'hff;
		rom[56]   	<= 8'hff;
		rom[57]   	<= 8'hff;
		rom[58]   	<= 8'hff;
		rom[59]   	<= 8'hff;
		rom[60]   	<= 8'hff;
		rom[61]   	<= 8'hff;
		rom[62]   	<= 8'hff;
		rom[63]   	<= 8'hff;
		rom[64]   	<= 8'hff;
		rom[65]   	<= 8'hff;
		rom[66]   	<= 8'hff;
		rom[67]   	<= 8'hff;
		rom[68]   	<= 8'hff;
		rom[69]   	<= 8'hff;
		rom[70]   	<= 8'hff;
		rom[71]   	<= 8'hff;
		rom[72]   	<= 8'hff;
		rom[73]   	<= 8'hff;
		rom[74]   	<= 8'hff;
		rom[75]   	<= 8'hff;
		rom[76]   	<= 8'hff;
		rom[77]   	<= 8'hff;
		rom[78]   	<= 8'hff;
		rom[79]   	<= 8'hff;
		rom[80]   	<= 8'hff;
		rom[81]   	<= 8'hff;
		rom[82]   	<= 8'hff;
		rom[83]   	<= 8'hff;
		rom[84]   	<= 8'hff;
		rom[85]   	<= 8'hff;
		rom[86]   	<= 8'hff;
		rom[87]   	<= 8'hff;
		rom[88]   	<= 8'hff;
		rom[89]   	<= 8'hff;
		rom[90]   	<= 8'hff;
		rom[91]   	<= 8'hff;
		rom[92]   	<= 8'hff;
		rom[93]   	<= 8'hff;
		rom[94]   	<= 8'hff;
		rom[95]   	<= 8'hff;
		rom[96]   	<= 8'hff;
		rom[97]   	<= 8'hff;
		rom[98]   	<= 8'hff;
		rom[99]   	<= 8'hff;
		rom[100]   	<= 8'hff;
		rom[101]   	<= 8'hff;
		rom[102]   	<= 8'hff;
		rom[103]   	<= 8'hff;
		rom[104]   	<= 8'hff;
		rom[105]   	<= 8'hff;
		rom[106]   	<= 8'hff;
		rom[107]   	<= 8'hff;
		rom[108]   	<= 8'hff;
		rom[109]   	<= 8'hff;
		rom[110]   	<= 8'hff;
		rom[111]   	<= 8'hff;
		rom[112]   	<= 8'hff;
		rom[113]   	<= 8'hff;
		rom[114]   	<= 8'hff;
		rom[115]   	<= 8'hff;
		rom[116]   	<= 8'hff;
		rom[117]   	<= 8'hff;
		rom[118]   	<= 8'hff;
		rom[119]   	<= 8'hff;
		rom[120]   	<= 8'hff;
		rom[121]   	<= 8'hff;
		rom[122]   	<= 8'hff;
		rom[123]   	<= 8'hff;
		rom[124]   	<= 8'hff;
		rom[125]   	<= 8'hff;
		rom[126]   	<= 8'hff;
		rom[127]   	<= 8'hff;
		rom[128]   	<= 8'hff;
		rom[129]   	<= 8'hff;
		rom[130]   	<= 8'hff;
		rom[131]   	<= 8'hff;
		rom[132]   	<= 8'hff;
		rom[133]   	<= 8'hff;
		rom[134]   	<= 8'hff;
		rom[135]   	<= 8'hff;
		rom[136]   	<= 8'hff;
		rom[137]   	<= 8'hff;
		rom[138]   	<= 8'hff;
		rom[139]   	<= 8'hff;
		rom[140]   	<= 8'hff;
		rom[141]   	<= 8'hff;
		rom[142]   	<= 8'hff;
		rom[143]   	<= 8'hff;
		rom[144]   	<= 8'hff;
		rom[145]   	<= 8'hff;
		rom[146]   	<= 8'hff;
		rom[147]   	<= 8'hff;
		rom[148]   	<= 8'hff;
		rom[149]   	<= 8'hff;
		rom[150]   	<= 8'hff;
		rom[151]   	<= 8'hff;
		rom[152]   	<= 8'hff;
		rom[153]   	<= 8'hff;
		rom[154]   	<= 8'hff;
		rom[155]   	<= 8'hff;
		rom[156]   	<= 8'hff;
		rom[157]   	<= 8'hff;
		rom[158]   	<= 8'hff;
		rom[159]   	<= 8'hff;
		rom[160]   	<= 8'hff;
		rom[161]   	<= 8'hff;
		rom[162]   	<= 8'hff;
		rom[163]   	<= 8'hff;
		rom[164]   	<= 8'hff;
		rom[165]   	<= 8'hff;
		rom[166]   	<= 8'hff;
		rom[167]   	<= 8'hff;
		rom[168]   	<= 8'hff;
		rom[169]   	<= 8'hff;
		rom[170]   	<= 8'hff;
		rom[171]   	<= 8'hff;
		rom[172]   	<= 8'hff;
		rom[173]   	<= 8'hff;
		rom[174]   	<= 8'hff;
		rom[175]   	<= 8'hff;
		rom[176]   	<= 8'hff;
		rom[177]   	<= 8'hff;
		rom[178]   	<= 8'hff;
		rom[179]   	<= 8'hff;
		rom[180]   	<= 8'hff;
		rom[181]   	<= 8'hff;
		rom[182]   	<= 8'hff;
		rom[183]   	<= 8'hff;
		rom[184]   	<= 8'hff;
		rom[185]   	<= 8'hff;
		rom[186]   	<= 8'hff;
		rom[187]   	<= 8'hff;
		rom[188]   	<= 8'hff;
		rom[189]   	<= 8'hff;
		rom[190]   	<= 8'hff;
		rom[191]   	<= 8'hff;
		rom[192]   	<= 8'hff;
		rom[193]   	<= 8'hff;
		rom[194]   	<= 8'hff;
		rom[195]   	<= 8'hff;
		rom[196]   	<= 8'hff;
		rom[197]   	<= 8'hff;
		rom[198]   	<= 8'hff;
		rom[199]   	<= 8'hff;
		rom[200]   	<= 8'hff;
		rom[201]   	<= 8'hff;
		rom[202]   	<= 8'hff;
		rom[203]   	<= 8'hff;
		rom[204]   	<= 8'hff;
		rom[205]   	<= 8'hff;
		rom[206]   	<= 8'hff;
		rom[207]   	<= 8'hff;
		rom[208]   	<= 8'hff;
		rom[209]   	<= 8'hff;
		rom[210]   	<= 8'hff;
		rom[211]   	<= 8'hff;
		rom[212]   	<= 8'hff;
		rom[213]   	<= 8'hff;
		rom[214]   	<= 8'hff;
		rom[215]   	<= 8'hff;
		rom[216]   	<= 8'hff;
		rom[217]   	<= 8'hff;
		rom[218]   	<= 8'hff;
		rom[219]   	<= 8'hff;
		rom[220]   	<= 8'hff;
		rom[221]   	<= 8'hff;
		rom[222]   	<= 8'hff;
		rom[223]   	<= 8'hff;
		rom[224]   	<= 8'hff;
		rom[225]   	<= 8'hff;
		rom[226]   	<= 8'hff;
		rom[227]   	<= 8'hff;
		rom[228]   	<= 8'hff;
		rom[229]   	<= 8'hff;
		rom[230]   	<= 8'hff;
		rom[231]   	<= 8'hff;
		rom[232]   	<= 8'hff;
		rom[233]   	<= 8'hff;
		rom[234]   	<= 8'hff;
		rom[235]   	<= 8'hff;
		rom[236]   	<= 8'hff;
		rom[237]   	<= 8'hff;
		rom[238]   	<= 8'hff;
		rom[239]   	<= 8'hff;
		rom[240]   	<= 8'hff;
		rom[241]   	<= 8'hff;
		rom[242]   	<= 8'hff;
		rom[243]   	<= 8'hff;
		rom[244]   	<= 8'hff;
		rom[245]   	<= 8'hff;
		rom[246]   	<= 8'hff;
		rom[247]   	<= 8'hff;
		rom[248]   	<= 8'hff;
		rom[249]   	<= 8'hff;
		rom[250]   	<= 8'hff;
		rom[251]   	<= 8'hff;
		rom[252]   	<= 8'hff;
		rom[253]   	<= 8'hff;
		rom[254]   	<= 8'hff;
		rom[255]   	<= 8'hff;
		rom[256]   	<= 8'hff;
		rom[257]   	<= 8'hff;
		rom[258]   	<= 8'hff;
		rom[259]   	<= 8'hff;
		rom[260]   	<= 8'hff;
		rom[261]   	<= 8'hff;
		rom[262]   	<= 8'hff;
		rom[263]   	<= 8'hff;
		rom[264]   	<= 8'hff;
		rom[265]   	<= 8'hff;
		rom[266]   	<= 8'hff;
		rom[267]   	<= 8'hff;
		rom[268]   	<= 8'hff;
		rom[269]   	<= 8'hff;
		rom[270]   	<= 8'hff;
		rom[271]   	<= 8'hff;
		rom[272]   	<= 8'hff;
		rom[273]   	<= 8'hff;
		rom[274]   	<= 8'hff;
		rom[275]   	<= 8'hff;
		rom[276]   	<= 8'hff;
		rom[277]   	<= 8'hff;
		rom[278]   	<= 8'hff;
		rom[279]   	<= 8'hff;
		rom[280]   	<= 8'hff;
		rom[281]   	<= 8'hff;
		rom[282]   	<= 8'hff;
		rom[283]   	<= 8'hff;
		rom[284]   	<= 8'hff;
		rom[285]   	<= 8'hff;
		rom[286]   	<= 8'hff;
		rom[287]   	<= 8'hff;
		rom[288]   	<= 8'hff;
		rom[289]   	<= 8'hff;
		rom[290]   	<= 8'hff;
		rom[291]   	<= 8'hff;
		rom[292]   	<= 8'hff;
		rom[293]   	<= 8'hff;
		rom[294]   	<= 8'hff;
		rom[295]   	<= 8'hff;
		rom[296]   	<= 8'hff;
		rom[297]   	<= 8'hff;
		rom[298]   	<= 8'hff;
		rom[299]   	<= 8'hff;
		rom[300]   	<= 8'hff;
		rom[301]   	<= 8'hff;
		rom[302]   	<= 8'hff;
		rom[303]   	<= 8'hff;
		rom[304]   	<= 8'hff;
		rom[305]   	<= 8'hff;
		rom[306]   	<= 8'hff;
		rom[307]   	<= 8'hff;
		rom[308]   	<= 8'hff;
		rom[309]   	<= 8'hff;
		rom[310]   	<= 8'hff;
		rom[311]   	<= 8'hff;
		rom[312]   	<= 8'hff;
		rom[313]   	<= 8'hff;
		rom[314]   	<= 8'hff;
		rom[315]   	<= 8'hff;
		rom[316]   	<= 8'hff;
		rom[317]   	<= 8'hff;
		rom[318]   	<= 8'hff;
		rom[319]   	<= 8'hff;
		rom[320]   	<= 8'hff;
		rom[321]   	<= 8'hff;
		rom[322]   	<= 8'hff;
		rom[323]   	<= 8'hff;
		rom[324]   	<= 8'hff;
		rom[325]   	<= 8'hff;
		rom[326]   	<= 8'hff;
		rom[327]   	<= 8'hff;
		rom[328]   	<= 8'hff;
		rom[329]   	<= 8'hff;
		rom[330]   	<= 8'hff;
		rom[331]   	<= 8'hff;
		rom[332]   	<= 8'hff;
		rom[333]   	<= 8'hff;
		rom[334]   	<= 8'hff;
		rom[335]   	<= 8'hff;
		rom[336]   	<= 8'hff;
		rom[337]   	<= 8'hff;
		rom[338]   	<= 8'hff;
		rom[339]   	<= 8'hff;
		rom[340]   	<= 8'hff;
		rom[341]   	<= 8'hff;
		rom[342]   	<= 8'hff;
		rom[343]   	<= 8'hff;
		rom[344]   	<= 8'hff;
		rom[345]   	<= 8'hff;
		rom[346]   	<= 8'hff;
		rom[347]   	<= 8'hff;
		rom[348]   	<= 8'hff;
		rom[349]   	<= 8'hff;
		rom[350]   	<= 8'hff;
		rom[351]   	<= 8'hff;
		rom[352]   	<= 8'hff;
		rom[353]   	<= 8'hff;
		rom[354]   	<= 8'hff;
		rom[355]   	<= 8'hff;
		rom[356]   	<= 8'hff;
		rom[357]   	<= 8'hff;
		rom[358]   	<= 8'hff;
		rom[359]   	<= 8'hff;
		rom[360]   	<= 8'hff;
		rom[361]   	<= 8'hff;
		rom[362]   	<= 8'hff;
		rom[363]   	<= 8'hff;
		rom[364]   	<= 8'hff;
		rom[365]   	<= 8'hff;
		rom[366]   	<= 8'hff;
		rom[367]   	<= 8'hff;
		rom[368]   	<= 8'hff;
		rom[369]   	<= 8'hff;
		rom[370]   	<= 8'hff;
		rom[371]   	<= 8'hff;
		rom[372]   	<= 8'hff;
		rom[373]   	<= 8'hff;
		rom[374]   	<= 8'hff;
		rom[375]   	<= 8'hff;
		rom[376]   	<= 8'hff;
		rom[377]   	<= 8'hff;
		rom[378]   	<= 8'hff;
		rom[379]   	<= 8'hff;
		rom[380]   	<= 8'hff;
		rom[381]   	<= 8'hff;
		rom[382]   	<= 8'hff;
		rom[383]   	<= 8'hff;
		rom[384]   	<= 8'hff;
		rom[385]   	<= 8'hff;
		rom[386]   	<= 8'hff;
		rom[387]   	<= 8'hff;
		rom[388]   	<= 8'hff;
		rom[389]   	<= 8'hff;
		rom[390]   	<= 8'hff;
		rom[391]   	<= 8'hff;
		rom[392]   	<= 8'hff;
		rom[393]   	<= 8'hff;
		rom[394]   	<= 8'hff;
		rom[395]   	<= 8'hff;
		rom[396]   	<= 8'hff;
		rom[397]   	<= 8'hff;
		rom[398]   	<= 8'hff;
		rom[399]   	<= 8'hff;
		rom[400]   	<= 8'hff;
		rom[401]   	<= 8'hff;
		rom[402]   	<= 8'hff;
		rom[403]   	<= 8'hff;
		rom[404]   	<= 8'hff;
		rom[405]   	<= 8'hff;
		rom[406]   	<= 8'hff;
		rom[407]   	<= 8'hff;
		rom[408]   	<= 8'hff;
		rom[409]   	<= 8'hff;
		rom[410]   	<= 8'hff;
		rom[411]   	<= 8'hff;
		rom[412]   	<= 8'hff;
		rom[413]   	<= 8'hff;
		rom[414]   	<= 8'hff;
		rom[415]   	<= 8'hff;
		rom[416]   	<= 8'hff;
		rom[417]   	<= 8'hff;
		rom[418]   	<= 8'hff;
		rom[419]   	<= 8'hff;
		rom[420]   	<= 8'hff;
		rom[421]   	<= 8'hff;
		rom[422]   	<= 8'hff;
		rom[423]   	<= 8'hff;
		rom[424]   	<= 8'hff;
		rom[425]   	<= 8'hff;
		rom[426]   	<= 8'hff;
		rom[427]   	<= 8'hff;
		rom[428]   	<= 8'hff;
		rom[429]   	<= 8'hff;
		rom[430]   	<= 8'hff;
		rom[431]   	<= 8'hff;
		rom[432]   	<= 8'hff;
		rom[433]   	<= 8'hff;
		rom[434]   	<= 8'hff;
		rom[435]   	<= 8'hff;
		rom[436]   	<= 8'hff;
		rom[437]   	<= 8'hff;
		rom[438]   	<= 8'hff;
		rom[439]   	<= 8'hff;
		rom[440]   	<= 8'hff;
		rom[441]   	<= 8'hff;
		rom[442]   	<= 8'hff;
		rom[443]   	<= 8'hff;
		rom[444]   	<= 8'hff;
		rom[445]   	<= 8'hff;
		rom[446]   	<= 8'hff;
		rom[447]   	<= 8'hff;
		rom[448]   	<= 8'hff;
		rom[449]   	<= 8'hff;
		rom[450]   	<= 8'hff;
		rom[451]   	<= 8'hff;
		rom[452]   	<= 8'hff;
		rom[453]   	<= 8'hff;
		rom[454]   	<= 8'hff;
		rom[455]   	<= 8'hff;
		rom[456]   	<= 8'hff;
		rom[457]   	<= 8'hff;
		rom[458]   	<= 8'hff;
		rom[459]   	<= 8'hff;
		rom[460]   	<= 8'hff;
		rom[461]   	<= 8'hff;
		rom[462]   	<= 8'hff;
		rom[463]   	<= 8'hff;
		rom[464]   	<= 8'hff;
		rom[465]   	<= 8'hff;
		rom[466]   	<= 8'hff;
		rom[467]   	<= 8'hff;
		rom[468]   	<= 8'hff;
		rom[469]   	<= 8'hff;
		rom[470]   	<= 8'hff;
		rom[471]   	<= 8'hff;
		rom[472]   	<= 8'hff;
		rom[473]   	<= 8'hff;
		rom[474]   	<= 8'hff;
		rom[475]   	<= 8'hff;
		rom[476]   	<= 8'hff;
		rom[477]   	<= 8'hff;
		rom[478]   	<= 8'hff;
		rom[479]   	<= 8'hff;
		rom[480]   	<= 8'hff;
		rom[481]   	<= 8'hff;
		rom[482]   	<= 8'hff;
		rom[483]   	<= 8'hff;
		rom[484]   	<= 8'hff;
		rom[485]   	<= 8'hff;
		rom[486]   	<= 8'hff;
		rom[487]   	<= 8'hff;
		rom[488]   	<= 8'hff;
		rom[489]   	<= 8'hff;
		rom[490]   	<= 8'hff;
		rom[491]   	<= 8'hff;
		rom[492]   	<= 8'hff;
		rom[493]   	<= 8'hff;
		rom[494]   	<= 8'hff;
		rom[495]   	<= 8'hff;
		rom[496]   	<= 8'hff;
		rom[497]   	<= 8'hff;
		rom[498]   	<= 8'hff;
		rom[499]   	<= 8'hff;
		rom[500]   	<= 8'hff;
		rom[501]   	<= 8'hff;
		rom[502]   	<= 8'hff;
		rom[503]   	<= 8'hff;
		rom[504]   	<= 8'hff;
		rom[505]   	<= 8'hff;
		rom[506]   	<= 8'hff;
		rom[507]   	<= 8'hff;
		rom[508]   	<= 8'hff;
		rom[509]   	<= 8'hff;
		rom[510]   	<= 8'hff;
		rom[511]   	<= 8'hff;
		rom[512]   	<= 8'hff;
		rom[513]   	<= 8'hff;
		rom[514]   	<= 8'hff;
		rom[515]   	<= 8'hff;
		rom[516]   	<= 8'hff;
		rom[517]   	<= 8'hff;
		rom[518]   	<= 8'hff;
		rom[519]   	<= 8'hff;
		rom[520]   	<= 8'hff;
		rom[521]   	<= 8'hff;
		rom[522]   	<= 8'hff;
		rom[523]   	<= 8'hff;
		rom[524]   	<= 8'hff;
		rom[525]   	<= 8'hff;
		rom[526]   	<= 8'hff;
		rom[527]   	<= 8'hff;
		rom[528]   	<= 8'hff;
		rom[529]   	<= 8'hff;
		rom[530]   	<= 8'hff;
		rom[531]   	<= 8'hff;
		rom[532]   	<= 8'hff;
		rom[533]   	<= 8'hff;
		rom[534]   	<= 8'hff;
		rom[535]   	<= 8'hff;
		rom[536]   	<= 8'hff;
		rom[537]   	<= 8'hff;
		rom[538]   	<= 8'hff;
		rom[539]   	<= 8'hff;
		rom[540]   	<= 8'hff;
		rom[541]   	<= 8'hff;
		rom[542]   	<= 8'hff;
		rom[543]   	<= 8'hff;
		rom[544]   	<= 8'hff;
		rom[545]   	<= 8'hff;
		rom[546]   	<= 8'hff;
		rom[547]   	<= 8'hff;
		rom[548]   	<= 8'hff;
		rom[549]   	<= 8'hff;
		rom[550]   	<= 8'hff;
		rom[551]   	<= 8'hff;
		rom[552]   	<= 8'hff;
		rom[553]   	<= 8'hff;
		rom[554]   	<= 8'hff;
		rom[555]   	<= 8'hff;
		rom[556]   	<= 8'hff;
		rom[557]   	<= 8'hff;
		rom[558]   	<= 8'hff;
		rom[559]   	<= 8'hff;
		rom[560]   	<= 8'hff;
		rom[561]   	<= 8'hff;
		rom[562]   	<= 8'hff;
		rom[563]   	<= 8'hff;
		rom[564]   	<= 8'hff;
		rom[565]   	<= 8'hff;
		rom[566]   	<= 8'hff;
		rom[567]   	<= 8'hff;
		rom[568]   	<= 8'hff;
		rom[569]   	<= 8'hff;
		rom[570]   	<= 8'hff;
		rom[571]   	<= 8'hff;
		rom[572]   	<= 8'hff;
		rom[573]   	<= 8'hff;
		rom[574]   	<= 8'hff;
		rom[575]   	<= 8'hff;
		rom[576]   	<= 8'hff;
		rom[577]   	<= 8'hff;
		rom[578]   	<= 8'hff;
		rom[579]   	<= 8'hff;
		rom[580]   	<= 8'hff;
		rom[581]   	<= 8'hff;
		rom[582]   	<= 8'hff;
		rom[583]   	<= 8'hff;
		rom[584]   	<= 8'hff;
		rom[585]   	<= 8'hff;
		rom[586]   	<= 8'hff;
		rom[587]   	<= 8'hff;
		rom[588]   	<= 8'hff;
		rom[589]   	<= 8'hff;
		rom[590]   	<= 8'hff;
		rom[591]   	<= 8'hff;
		rom[592]   	<= 8'hff;
		rom[593]   	<= 8'hff;
		rom[594]   	<= 8'hff;
		rom[595]   	<= 8'hff;
		rom[596]   	<= 8'hff;
		rom[597]   	<= 8'hff;
		rom[598]   	<= 8'hff;
		rom[599]   	<= 8'hff;
		rom[600]   	<= 8'hff;
		rom[601]   	<= 8'hff;
		rom[602]   	<= 8'hff;
		rom[603]   	<= 8'hff;
		rom[604]   	<= 8'hff;
		rom[605]   	<= 8'hff;
		rom[606]   	<= 8'hff;
		rom[607]   	<= 8'hff;
		rom[608]   	<= 8'hff;
		rom[609]   	<= 8'hff;
		rom[610]   	<= 8'hff;
		rom[611]   	<= 8'hff;
		rom[612]   	<= 8'hff;
		rom[613]   	<= 8'hff;
		rom[614]   	<= 8'hff;
		rom[615]   	<= 8'hff;
		rom[616]   	<= 8'hff;
		rom[617]   	<= 8'hff;
		rom[618]   	<= 8'hff;
		rom[619]   	<= 8'hff;
		rom[620]   	<= 8'hff;
		rom[621]   	<= 8'hff;
		rom[622]   	<= 8'hff;
		rom[623]   	<= 8'hff;
		rom[624]   	<= 8'hff;
		rom[625]   	<= 8'hff;
		rom[626]   	<= 8'hff;
		rom[627]   	<= 8'hff;
		rom[628]   	<= 8'hff;
		rom[629]   	<= 8'hff;
		rom[630]   	<= 8'hff;
		rom[631]   	<= 8'hff;
		rom[632]   	<= 8'hff;
		rom[633]   	<= 8'hff;
		rom[634]   	<= 8'hff;
		rom[635]   	<= 8'hff;
		rom[636]   	<= 8'hff;
		rom[637]   	<= 8'hff;
		rom[638]   	<= 8'hff;
		rom[639]   	<= 8'hff;
		rom[640]   	<= 8'hff;
		rom[641]   	<= 8'hff;
		rom[642]   	<= 8'hff;
		rom[643]   	<= 8'hff;
		rom[644]   	<= 8'hff;
		rom[645]   	<= 8'hff;
		rom[646]   	<= 8'hff;
		rom[647]   	<= 8'hff;
		rom[648]   	<= 8'hff;
		rom[649]   	<= 8'hff;
		rom[650]   	<= 8'hff;
		rom[651]   	<= 8'hff;
		rom[652]   	<= 8'hff;
		rom[653]   	<= 8'hff;
		rom[654]   	<= 8'hff;
		rom[655]   	<= 8'hff;
		rom[656]   	<= 8'hff;
		rom[657]   	<= 8'hff;
		rom[658]   	<= 8'hff;
		rom[659]   	<= 8'hff;
		rom[660]   	<= 8'hff;
		rom[661]   	<= 8'hff;
		rom[662]   	<= 8'hff;
		rom[663]   	<= 8'hff;
		rom[664]   	<= 8'hff;
		rom[665]   	<= 8'hff;
		rom[666]   	<= 8'hff;
		rom[667]   	<= 8'hff;
		rom[668]   	<= 8'hff;
		rom[669]   	<= 8'hff;
		rom[670]   	<= 8'hff;
		rom[671]   	<= 8'hff;
		rom[672]   	<= 8'hff;
		rom[673]   	<= 8'hff;
		rom[674]   	<= 8'hff;
		rom[675]   	<= 8'hff;
		rom[676]   	<= 8'hff;
		rom[677]   	<= 8'hff;
		rom[678]   	<= 8'hff;
		rom[679]   	<= 8'hff;
		rom[680]   	<= 8'hff;
		rom[681]   	<= 8'hff;
		rom[682]   	<= 8'hff;
		rom[683]   	<= 8'hff;
		rom[684]   	<= 8'hff;
		rom[685]   	<= 8'hff;
		rom[686]   	<= 8'hff;
		rom[687]   	<= 8'hff;
		rom[688]   	<= 8'hff;
		rom[689]   	<= 8'hff;
		rom[690]   	<= 8'hff;
		rom[691]   	<= 8'hff;
		rom[692]   	<= 8'hff;
		rom[693]   	<= 8'hff;
		rom[694]   	<= 8'hff;
		rom[695]   	<= 8'hff;
		rom[696]   	<= 8'hff;
		rom[697]   	<= 8'hff;
		rom[698]   	<= 8'hff;
		rom[699]   	<= 8'hff;
		rom[700]   	<= 8'hff;
		rom[701]   	<= 8'hff;
		rom[702]   	<= 8'hff;
		rom[703]   	<= 8'hff;
		rom[704]   	<= 8'hff;
		rom[705]   	<= 8'hff;
		rom[706]   	<= 8'hff;
		rom[707]   	<= 8'hff;
		rom[708]   	<= 8'hff;
		rom[709]   	<= 8'hff;
		rom[710]   	<= 8'hff;
		rom[711]   	<= 8'hff;
		rom[712]   	<= 8'hff;
		rom[713]   	<= 8'hff;
		rom[714]   	<= 8'hff;
		rom[715]   	<= 8'hff;
		rom[716]   	<= 8'hff;
		rom[717]   	<= 8'hff;
		rom[718]   	<= 8'hff;
		rom[719]   	<= 8'hff;
		rom[720]   	<= 8'hff;
		rom[721]   	<= 8'hff;
		rom[722]   	<= 8'hff;
		rom[723]   	<= 8'hff;
		rom[724]   	<= 8'hff;
		rom[725]   	<= 8'hff;
		rom[726]   	<= 8'hff;
		rom[727]   	<= 8'hff;
		rom[728]   	<= 8'hff;
		rom[729]   	<= 8'hff;
		rom[730]   	<= 8'hff;
		rom[731]   	<= 8'hff;
		rom[732]   	<= 8'hff;
		rom[733]   	<= 8'hff;
		rom[734]   	<= 8'hff;
		rom[735]   	<= 8'hff;
		rom[736]   	<= 8'hff;
		rom[737]   	<= 8'hff;
		rom[738]   	<= 8'hff;
		rom[739]   	<= 8'hff;
		rom[740]   	<= 8'hff;
		rom[741]   	<= 8'hff;
		rom[742]   	<= 8'hff;
		rom[743]   	<= 8'hff;
		rom[744]   	<= 8'hff;
		rom[745]   	<= 8'hff;
		rom[746]   	<= 8'hff;
		rom[747]   	<= 8'hff;
		rom[748]   	<= 8'hff;
		rom[749]   	<= 8'hff;
		rom[750]   	<= 8'hff;
		rom[751]   	<= 8'hff;
		rom[752]   	<= 8'hff;
		rom[753]   	<= 8'hff;
		rom[754]   	<= 8'hff;
		rom[755]   	<= 8'hff;
		rom[756]   	<= 8'hff;
		rom[757]   	<= 8'hff;
		rom[758]   	<= 8'hff;
		rom[759]   	<= 8'hff;
		rom[760]   	<= 8'hff;
		rom[761]   	<= 8'hff;
		rom[762]   	<= 8'hff;
		rom[763]   	<= 8'hff;
		rom[764]   	<= 8'hff;
		rom[765]   	<= 8'hff;
		rom[766]   	<= 8'hff;
		rom[767]   	<= 8'hff;
		rom[768]   	<= 8'hff;
		rom[769]   	<= 8'hff;
		rom[770]   	<= 8'hff;
		rom[771]   	<= 8'hff;
		rom[772]   	<= 8'hff;
		rom[773]   	<= 8'hff;
		rom[774]   	<= 8'hff;
		rom[775]   	<= 8'hff;
		rom[776]   	<= 8'hff;
		rom[777]   	<= 8'hff;
		rom[778]   	<= 8'hff;
		rom[779]   	<= 8'hff;
		rom[780]   	<= 8'hff;
		rom[781]   	<= 8'hff;
		rom[782]   	<= 8'hff;
		rom[783]   	<= 8'hff;
		rom[784]   	<= 8'hff;
		rom[785]   	<= 8'hff;
		rom[786]   	<= 8'hff;
		rom[787]   	<= 8'hff;
		rom[788]   	<= 8'hff;
		rom[789]   	<= 8'hff;
		rom[790]   	<= 8'hff;
		rom[791]   	<= 8'hff;
		rom[792]   	<= 8'hff;
		rom[793]   	<= 8'hff;
		rom[794]   	<= 8'hff;
		rom[795]   	<= 8'hff;
		rom[796]   	<= 8'hff;
		rom[797]   	<= 8'hff;
		rom[798]   	<= 8'hff;
		rom[799]   	<= 8'hff;
		rom[800]   	<= 8'hff;
		rom[801]   	<= 8'hff;
		rom[802]   	<= 8'hff;
		rom[803]   	<= 8'hff;
		rom[804]   	<= 8'hff;
		rom[805]   	<= 8'hff;
		rom[806]   	<= 8'hff;
		rom[807]   	<= 8'hff;
		rom[808]   	<= 8'hff;
		rom[809]   	<= 8'hff;
		rom[810]   	<= 8'hff;
		rom[811]   	<= 8'hff;
		rom[812]   	<= 8'hff;
		rom[813]   	<= 8'hff;
		rom[814]   	<= 8'hff;
		rom[815]   	<= 8'hff;
		rom[816]   	<= 8'hff;
		rom[817]   	<= 8'hff;
		rom[818]   	<= 8'hff;
		rom[819]   	<= 8'hff;
		rom[820]   	<= 8'hff;
		rom[821]   	<= 8'hff;
		rom[822]   	<= 8'hff;
		rom[823]   	<= 8'hff;
		rom[824]   	<= 8'hff;
		rom[825]   	<= 8'hff;
		rom[826]   	<= 8'hff;
		rom[827]   	<= 8'hff;
		rom[828]   	<= 8'hff;
		rom[829]   	<= 8'hff;
		rom[830]   	<= 8'hff;
		rom[831]   	<= 8'hff;
		rom[832]   	<= 8'hff;
		rom[833]   	<= 8'hff;
		rom[834]   	<= 8'hff;
		rom[835]   	<= 8'hff;
		rom[836]   	<= 8'hff;
		rom[837]   	<= 8'hff;
		rom[838]   	<= 8'hff;
		rom[839]   	<= 8'hff;
		rom[840]   	<= 8'hff;
		rom[841]   	<= 8'hff;
		rom[842]   	<= 8'hff;
		rom[843]   	<= 8'hff;
		rom[844]   	<= 8'hff;
		rom[845]   	<= 8'hff;
		rom[846]   	<= 8'hff;
		rom[847]   	<= 8'hff;
		rom[848]   	<= 8'hff;
		rom[849]   	<= 8'hff;
		rom[850]   	<= 8'hff;
		rom[851]   	<= 8'hff;
		rom[852]   	<= 8'hff;
		rom[853]   	<= 8'hff;
		rom[854]   	<= 8'hff;
		rom[855]   	<= 8'hff;
		rom[856]   	<= 8'hff;
		rom[857]   	<= 8'hff;
		rom[858]   	<= 8'hff;
		rom[859]   	<= 8'hff;
		rom[860]   	<= 8'hff;
		rom[861]   	<= 8'hff;
		rom[862]   	<= 8'hff;
		rom[863]   	<= 8'hff;
		rom[864]   	<= 8'hff;
		rom[865]   	<= 8'hff;
		rom[866]   	<= 8'hff;
		rom[867]   	<= 8'hff;
		rom[868]   	<= 8'hff;
		rom[869]   	<= 8'hff;
		rom[870]   	<= 8'hff;
		rom[871]   	<= 8'hff;
		rom[872]   	<= 8'hff;
		rom[873]   	<= 8'hff;
		rom[874]   	<= 8'hff;
		rom[875]   	<= 8'hff;
		rom[876]   	<= 8'hff;
		rom[877]   	<= 8'hff;
		rom[878]   	<= 8'hff;
		rom[879]   	<= 8'hff;
		rom[880]   	<= 8'hff;
		rom[881]   	<= 8'hff;
		rom[882]   	<= 8'hff;
		rom[883]   	<= 8'hff;
		rom[884]   	<= 8'hff;
		rom[885]   	<= 8'hff;
		rom[886]   	<= 8'hff;
		rom[887]   	<= 8'hff;
		rom[888]   	<= 8'hff;
		rom[889]   	<= 8'hff;
		rom[890]   	<= 8'hff;
		rom[891]   	<= 8'hff;
		rom[892]   	<= 8'hff;
		rom[893]   	<= 8'hff;
		rom[894]   	<= 8'hff;
		rom[895]   	<= 8'hff;
		rom[896]   	<= 8'hff;
		rom[897]   	<= 8'hff;
		rom[898]   	<= 8'hff;
		rom[899]   	<= 8'hff;
		rom[900]   	<= 8'hff;
		rom[901]   	<= 8'hff;
		rom[902]   	<= 8'hff;
		rom[903]   	<= 8'hff;
		rom[904]   	<= 8'hff;
		rom[905]   	<= 8'hff;
		rom[906]   	<= 8'hff;
		rom[907]   	<= 8'hff;
		rom[908]   	<= 8'hff;
		rom[909]   	<= 8'hff;
		rom[910]   	<= 8'hff;
		rom[911]   	<= 8'hff;
		rom[912]   	<= 8'hff;
		rom[913]   	<= 8'hff;
		rom[914]   	<= 8'hff;
		rom[915]   	<= 8'hff;
		rom[916]   	<= 8'hff;
		rom[917]   	<= 8'hff;
		rom[918]   	<= 8'hff;
		rom[919]   	<= 8'hff;
		rom[920]   	<= 8'hff;
		rom[921]   	<= 8'hff;
		rom[922]   	<= 8'hff;
		rom[923]   	<= 8'hff;
		rom[924]   	<= 8'hff;
		rom[925]   	<= 8'hff;
		rom[926]   	<= 8'hff;
		rom[927]   	<= 8'hff;
		rom[928]   	<= 8'hff;
		rom[929]   	<= 8'hff;
		rom[930]   	<= 8'hff;
		rom[931]   	<= 8'hff;
		rom[932]   	<= 8'hff;
		rom[933]   	<= 8'hff;
		rom[934]   	<= 8'hff;
		rom[935]   	<= 8'hff;
		rom[936]   	<= 8'hff;
		rom[937]   	<= 8'hff;
		rom[938]   	<= 8'hff;
		rom[939]   	<= 8'hff;
		rom[940]   	<= 8'hff;
		rom[941]   	<= 8'hff;
		rom[942]   	<= 8'hff;
		rom[943]   	<= 8'hff;
		rom[944]   	<= 8'hff;
		rom[945]   	<= 8'hff;
		rom[946]   	<= 8'hff;
		rom[947]   	<= 8'hff;
		rom[948]   	<= 8'hff;
		rom[949]   	<= 8'hff;
		rom[950]   	<= 8'hff;
		rom[951]   	<= 8'hff;
		rom[952]   	<= 8'hff;
		rom[953]   	<= 8'hff;
		rom[954]   	<= 8'hff;
		rom[955]   	<= 8'hff;
		rom[956]   	<= 8'hff;
		rom[957]   	<= 8'hff;
		rom[958]   	<= 8'hff;
		rom[959]   	<= 8'hff;
		rom[960]   	<= 8'hff;
		rom[961]   	<= 8'hff;
		rom[962]   	<= 8'hff;
		rom[963]   	<= 8'hff;
		rom[964]   	<= 8'hff;
		rom[965]   	<= 8'hff;
		rom[966]   	<= 8'hff;
		rom[967]   	<= 8'hff;
		rom[968]   	<= 8'hff;
		rom[969]   	<= 8'hff;
		rom[970]   	<= 8'hff;
		rom[971]   	<= 8'hff;
		rom[972]   	<= 8'hff;
		rom[973]   	<= 8'hff;
		rom[974]   	<= 8'hff;
		rom[975]   	<= 8'hff;
		rom[976]   	<= 8'hff;
		rom[977]   	<= 8'hff;
		rom[978]   	<= 8'hff;
		rom[979]   	<= 8'hff;
		rom[980]   	<= 8'hff;
		rom[981]   	<= 8'hff;
		rom[982]   	<= 8'hff;
		rom[983]   	<= 8'hff;
		rom[984]   	<= 8'hff;
		rom[985]   	<= 8'hff;
		rom[986]   	<= 8'hff;
		rom[987]   	<= 8'hff;
		rom[988]   	<= 8'hff;
		rom[989]   	<= 8'hff;
		rom[990]   	<= 8'hff;
		rom[991]   	<= 8'hff;
		rom[992]   	<= 8'hff;
		rom[993]   	<= 8'hff;
		rom[994]   	<= 8'hff;
		rom[995]   	<= 8'hff;
		rom[996]   	<= 8'hff;
		rom[997]   	<= 8'hff;
		rom[998]   	<= 8'hff;
		rom[999]   	<= 8'hff;
		rom[1000]	<= 8'hff;
		rom[1001]	<= 8'hff;
		rom[1002]	<= 8'hff;
		rom[1003]	<= 8'hff;
		rom[1004]	<= 8'hff;
		rom[1005]	<= 8'hff;
		rom[1006]	<= 8'hff;
		rom[1007]	<= 8'hff;
		rom[1008]	<= 8'hff;
		rom[1009]	<= 8'hff;
		rom[1010]	<= 8'hff;
		rom[1011]	<= 8'hff;
		rom[1012]	<= 8'hff;
		rom[1013]	<= 8'hff;
		rom[1014]	<= 8'hff;
		rom[1015]	<= 8'hff;
		rom[1016]	<= 8'hff;
		rom[1017]	<= 8'hff;
		rom[1018]	<= 8'hff;
		rom[1019]	<= 8'hff;
		rom[1020]	<= 8'hff;
		rom[1021]	<= 8'hff;
		rom[1022]	<= 8'hff;
		rom[1023]	<= 8'hff;
end

endmodule
